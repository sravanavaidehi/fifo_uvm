class f_sqr extends uvm_sequencer #(item);
  `uvm_component_utils(f_sqr)
  function new(string name = "f_sqr", uvm_component parent = null);
    super.new(name,parent);
  endfunction
endclass

            
